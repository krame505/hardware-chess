package Driver where

import Chess
import SearchCore
import GenCMsg
import GenCRepr
import GetPut
import ClientServer
import Connectable
import COBS
import CShow

data Command = GetState
             | Move Move
             | GetSearchMove { rid :: RequestId; depth :: Depth; }
             | CancelSearch
             | Reset
  deriving (Bits)

interface ChessMsgs =
  command :: Rx 2 2 Command
  state :: Tx 2 2 State
  outcome :: Tx 2 2 Outcome
  moves :: Tx 64 8 MoveResponse
  searchResult :: Tx 2 2 SearchResult

interface ChessDriver =
  txData :: Get (Bit 8)
  rxData :: Put (Bit 8)

  status :: Bit 16  {-# always_ready, always_enabled #-}

{-# verilog mkChessDriver #-}
mkChessDriver :: Module ChessDriver
mkChessDriver = _mkChessDriver

-- Seperate due to the context
_mkChessDriver :: (GenCMsg ChessMsgs rxBytes txBytes) => Module ChessDriver
_mkChessDriver = module
  writeCMsgDecls "chess" (_ :: ChessMsgs)

  enc :: COBSEncoder txBytes <- mkCOBSEncoder
  dec :: COBSDecoder rxBytes <- mkCOBSDecoder
  msgMgr :: MsgManager ChessMsgs rxBytes txBytes <- mkMsgManager

  dec.msg <-> dropSize msgMgr.rxMsg
  msgMgr.txMsg <-> enc.msg

  state :: Reg State <- mkReg initialState
  moveUpdate <- mkMoveUpdate
  searchCore <- mkParallelSearchCore

  searchCore.moves <-> toPut msgMgr.fifos.moves

  let updateState newState = do
        state := newState
        searchCore.server.request.put $ defaultValue {rid=0; state=newState; depth=1; getMoves=True;}
        msgMgr.fifos.state.enq newState

      commandRules =
        rules
          "handle_GetState": when GetState <- msgMgr.fifos.command.first ==> do
            $display "handle_GetState"
            updateState state
            msgMgr.fifos.command.deq
          "handle_Move": when Move m <- msgMgr.fifos.command.first ==> do
            $display "handle_Move"
            moveUpdate.enq state m
            msgMgr.fifos.command.deq
          "handle_GetSearchMove": when GetSearchMove {rid=rid; depth=depth;} <- msgMgr.fifos.command.first ==> do
            $display "handle_GetSearchMove"
            searchCore.server.request.put $ defaultValue {rid=rid; state=state; depth=depth;}
            msgMgr.fifos.command.deq
          "handle_CancelSearch": when CancelSearch <- msgMgr.fifos.command.first ==> do
            $display "handle_CancelSearch"
            searchCore.clear
            msgMgr.fifos.command.deq
          "handle_Reset": when Reset <- msgMgr.fifos.command.first ==> do
            $display "handle_Reset"
            updateState $ initialState
            msgMgr.fifos.command.deq

      updateRules =
        rules
          "report_move_update": when True ==> do
            $display "report_move_update"
            updateState moveUpdate.nextState
            moveUpdate.deq

          "report_search_outcome": when True ==> do
            $display "report_search_outcome"
            result <- searchCore.server.response.get
            if result.rid == 0
              then msgMgr.fifos.outcome.enq result.outcome
              else msgMgr.fifos.searchResult.enq result

  addRules $ commandRules `rJoinDescendingUrgency` updateRules

  interface
    txData = enc.byte
    rxData = dec.byte
    status = searchCore.status
