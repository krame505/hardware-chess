package Driver where

import Chess
import GenCMsg
import GenCRepr
import GetPut
import Connectable
import COBS
import CShow

data Command = GetState
             | Move Move
             | Reset
  deriving (Bits)

interface ChessMsgs =
  command :: Rx 2 2 Command
  state :: Tx 2 2 State
  moves :: Tx 64 8 MoveResponse

interface ChessDriver =
  txData :: Get (Bit 8)
  rxData :: Put (Bit 8)

mkChessDriver :: (GenCMsg ChessMsgs rxBytes txBytes) => Module ChessDriver
mkChessDriver = module
  writeCMsgDecls "chess" (_ :: ChessMsgs)

  enc :: COBSEncoder txBytes <- mkCOBSEncoder
  dec :: COBSDecoder rxBytes <- mkCOBSDecoder
  msgMgr :: MsgManager ChessMsgs rxBytes txBytes <- mkMsgManager

  dec.msg <-> dropSize msgMgr.rxMsg
  msgMgr.txMsg <-> enc.msg

  state :: Reg State <- mkReg initialState
  stateUpdate :: RWire State <- mkRWire

  eval :: StateEval <- mkStateEval
  eval.moves <-> toPut msgMgr.fifos.moves

  rules
    "handle_GetState": when GetState <- msgMgr.fifos.command.first ==> do
      stateUpdate.wset state
      msgMgr.fifos.command.deq
    "handle_Move": when Move m <- msgMgr.fifos.command.first ==> do
      stateUpdate.wset $ move m state
      msgMgr.fifos.command.deq
    "handle_Reset": when Reset <- msgMgr.fifos.command.first ==> do
      stateUpdate.wset initialState
      msgMgr.fifos.command.deq
    "update_state": when Just newState <- stateUpdate.wget ==> do
      state := newState
      eval.state.put newState
      msgMgr.fifos.state.enq newState

  interface
    txData = enc.byte
    rxData = dec.byte
