package HwTop where

import Driver
import RS232
import GetPut
import Connectable
import Clocks

interface Top =
  tx :: Bit 1 {-# always_ready, always_enabled #-}
  rx :: Bit 1 -> Action {-# always_ready, always_enabled, prefix="", arg_names = [rx] #-}
  status :: Bit 8 {-# always_ready, always_enabled #-}

clockFreq :: Integer
clockFreq = 100000000

clockDivisor :: Integer
clockDivisor = 5

baud :: Integer
baud = 115200

{-# verilog mkTop #-}
mkTop :: Module Top
mkTop = module
  clockDivider <- mkClockDivider clockDivisor
  reset <- mkReset clockDivisor True clockDivider.slowClock
  driver <- changeSpecialWires (Just clockDivider.slowClock) (Just reset.new_rst) Nothing mkChessDriver
  driverTx <- mkConverter 2 driver.txData
  driverRx <- mkConverter 2 driver.rxData

  uart :: UART 8 <- mkUART 8 NONE STOP_1 (fromInteger $ clockFreq / (baud * 16))

  -- Wait for first byte to be recieved before sending data
  writeEnable <- mkReg False
  rules
    "tx": when writeEnable ==> do
      c <- driverTx.get
      uart.rx.put c

    "rx": when True ==> do
      c <- uart.tx.get
      driverRx.put $ truncate $ pack c
      writeEnable := True

  driverStatus <- mkConverter 2 $ toGet driver.status
  lastStatus :: Reg (Bit 8) <- mkReg 0
  driverStatus <-> toPut lastStatus._write

  interface
    tx = uart.rs232.sout
    rx = uart.rs232.sin
    status = lastStatus
