package SearchCore where

import Chess
import FIFO
import FIFOF
import BRAMFIFO
import GetPut
import Connectable
import Vector
import CShow

type Depth = UInt 8
type Score = Int 8
type MoveCount = UInt 8

padDepth :: Depth -> String
padDepth 10 = "                    "
padDepth 9 = "                  "
padDepth 8 = "                "
padDepth 7 = "              "
padDepth 6 = "            "
padDepth 5 = "          "
padDepth 4 = "        "
padDepth 3 = "      "
padDepth 2 = "    "
padDepth 1 = "  "
padDepth _ = ""

pieceValue :: PieceKind -> Score
pieceValue Pawn = 1
pieceValue Knight = 3
pieceValue Bishop = 3
pieceValue Rook = 5
pieceValue Queen = 9
pieceValue King = 0

heuristicScore :: State -> Score
heuristicScore state =
  let squareScore Nothing = 0
      squareScore (Just piece) =
        (if piece.color == state.turn then id else negate) $ pieceValue piece.kind
  in foldr1 (+) $ map squareScore $ concat state.board

struct SearchQuery =
  state :: State
  depth :: Depth
 deriving (Bits)

struct SearchResult =
  bestMove :: Maybe Move
  score :: Score
  depth :: Depth
 deriving (Bits)

interface Frame =
  putState :: State -> Bool -> Action
  putScore :: Score -> ActionValue Bool
  state :: State
  hasMove :: Bool
  score :: Score
  moves :: FIFOF Move

mkFrame :: Module Frame
mkFrame = module
  state <- mkReg _
  inCheck <- mkReg False
  moves <- {- mkSizedBRAMFIFOF -} mkSizedFIFOF maxStateMoves
  hasMove <- mkReg False
  bestScore <- mkReg 0
  interface
    putState s c =
      do state := s
         inCheck := c
         hasMove := False
    putScore s =
      do hasMove := True
         let isBestScore = s > bestScore || not hasMove
         if isBestScore then bestScore := s else noAction
         return isBestScore
    state = state
    hasMove = hasMove
    score =
      if hasMove then bestScore
      else if inCheck then minBound + 1  -- Checkmate
      else 0  -- Draw
    moves = moves

interface (SearchCore :: # -> *) maxDepth =
  query :: Put SearchQuery
  result :: Get SearchResult

mkSearchCore :: Module (SearchCore maxDepth)
mkSearchCore = module
  queries :: FIFO SearchQuery <- mkFIFO
  results :: FIFO SearchResult <- mkFIFO

  initialDepth :: Reg Depth <- mkReg 0

  stack :: Vector maxDepth Frame <- replicateM mkFrame
  stackSize :: Reg Depth <- mkReg 0
  let depth = initialDepth - stackSize
      nextFrame = select stack stackSize
      topFrame = select stack (stackSize - 1)
      prevFrame = select stack (stackSize - 2)

  state :: Wire State <- mkWire
  stateHeuristicScore :: Wire Score <- mkWire
  currentPlayerInCheck :: Wire Bool <- mkWire
  otherPlayerInCheck :: Wire Bool <- mkWire

  eval :: MoveEval <- mkMoveEval
  movesComplete :: Reg Bool <- mkReg True
  let putState = do
        nextFrame.putState state otherPlayerInCheck
        eval.state.put state
        movesComplete := False

  bestMove :: Reg Move <- mkReg _
  currentMove :: Reg Move <- mkReg _

  rules
    "gen_state": when stackSize > 0 ==> state := move topFrame.moves.first topFrame.state
    "use_query_state": when stackSize == 0 ==> state := queries.first.state
    "eval_state": when True ==> do
      stateHeuristicScore := heuristicScore state
      currentPlayerInCheck := inCheck state.board topFrame.state.turn
      otherPlayerInCheck := inCheck state.board (otherColor topFrame.state.turn)

    "put_NextMove": when not movesComplete, NextMove m <- eval.move.first ==> do
      -- $display (padDepth stackSize) stackSize " put_NextMove " (cshow m)
      topFrame.moves.enq m
      eval.move.deq
    "put_NoMove": when not movesComplete, NoMove <- eval.move.first ==> do
      -- $display (padDepth stackSize) stackSize " put_NoMove"
      movesComplete := True
      eval.move.deq

    "ignore_check_state": when stackSize > 0, currentPlayerInCheck ==> do
      $display (padDepth stackSize) stackSize " ignore_check_state " (cshow topFrame.moves.first)
      topFrame.moves.deq

    "heuristic_state": when stackSize > 0, not currentPlayerInCheck, depth == 0 ==> do
      $display (padDepth stackSize) stackSize " heuristic_state " (cshow topFrame.moves.first) " " stateHeuristicScore
      topFrame.putScore $ negate stateHeuristicScore
      topFrame.moves.deq

    when movesComplete
      rules
        "push_state": when stackSize > 0, not currentPlayerInCheck, depth > 0 ==> do
          $display (padDepth stackSize) stackSize " push_state " (cshow topFrame.moves.first) " " stateHeuristicScore
          putState
          if stackSize == 1 then currentMove := topFrame.moves.first else noAction
          topFrame.moves.deq
          stackSize := stackSize + 1

        "pop_state": when stackSize > 1, not topFrame.moves.notEmpty ==> do
          $display (padDepth stackSize) stackSize " pop_state " topFrame.score
          isBestScore <- prevFrame.putScore $ negate topFrame.score
          if stackSize == 2 && isBestScore then bestMove := currentMove else noAction
          stackSize := stackSize - 1

        "push_query_state": when stackSize == 0 ==> do
          $display (padDepth stackSize) stackSize " push_query_state " (cshow queries.first)
          initialDepth := queries.first.depth
          putState
          stackSize := 1
          queries.deq

        "pop_result_state": when stackSize == 1, not topFrame.moves.notEmpty ==> do
          let result = SearchResult {
                bestMove = if topFrame.hasMove then Just bestMove else Nothing;
                score=topFrame.score;
                depth=initialDepth;
              }
          $display (padDepth stackSize) stackSize " pop_result_state " (cshow result)
          results.enq result
          stackSize := 0

  interface
    query = toPut queries
    result = toGet results

{-# verilog mkDefaultSearchCore #-}
mkDefaultSearchCore :: Module (SearchCore 3)
mkDefaultSearchCore = mkSearchCore
