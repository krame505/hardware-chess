package Driver where

import GetPut

interface Driver =
  txData :: Get (Bit 8)
  rxData :: Put (Bit 8)

  status :: Bit 16  {-# always_ready, always_enabled #-}
