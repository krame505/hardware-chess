package VSimTop where

import Chess
import SearchCore
import CShow
import GetPut
import ClientServer

searchDepth :: Depth
searchDepth = 3

{-# verilog sysChessVSim #-}
sysChessVSim :: Module Empty
sysChessVSim = module
  searchCore <- mkParallelSearchCore
  moveUpdate <- mkMoveUpdate
  state <- mkReg initialState

  init <- mkReg False
  rules
    "init": when not init ==> do
      $display (cshow state)
      searchCore.server.request.put $ SearchQuery {rid=0; state=state; depth=searchDepth; getMoves=False; alpha=Nothing; beta=Nothing;}
      init := True
    "get_result": when init ==> do
      result <- searchCore.server.response.get
      $display (cshow result)
      case result.bestMove of
        Just m -> do
          moveUpdate.putState state
          moveUpdate.putMove m
        Nothing -> $finish
    "put_query": when init ==> do
      $display moveUpdate.newState
      state := moveUpdate.newState
      searchCore.server.request.put $ SearchQuery {rid=0; state=moveUpdate.newState; depth=searchDepth; getMoves=False; alpha=Nothing; beta=Nothing;}
