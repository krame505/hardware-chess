package Driver where

import Chess
import SearchCore
import GenCMsg
import GenCRepr
import GetPut
import Connectable
import COBS
import CShow

searchDepth :: Depth
searchDepth = 3

data Command = GetState
             | Move Move
             | GetSearchMove
             | Reset
  deriving (Bits)

data Outcome = NoOutcome | Check | CheckMate | Draw
  deriving (Bits)

interface ChessMsgs =
  command :: Rx 2 2 Command
  state :: Tx 2 2 State
  outcome :: Tx 2 2 Outcome
  moves :: Tx 64 8 MoveResponse
  searchMove :: Tx 2 2 (Maybe Move)

interface ChessDriver =
  txData :: Get (Bit 8)
  rxData :: Put (Bit 8)

{-# verilog mkChessDriver #-}
mkChessDriver :: Module ChessDriver
mkChessDriver = _mkChessDriver

-- Seperate due to the context
_mkChessDriver :: (GenCMsg ChessMsgs rxBytes txBytes) => Module ChessDriver
_mkChessDriver = module
  writeCMsgDecls "chess" (_ :: ChessMsgs)

  enc :: COBSEncoder txBytes <- mkCOBSEncoder
  dec :: COBSDecoder rxBytes <- mkCOBSDecoder
  msgMgr :: MsgManager ChessMsgs rxBytes txBytes <- mkMsgManager

  dec.msg <-> dropSize msgMgr.rxMsg
  msgMgr.txMsg <-> enc.msg

  state :: Reg State <- mkReg initialState
  eval :: MoveEval <- mkMoveEval
  searchCore <- mkDefaultSearchCore
  let updateState newState = do
        state := newState
        eval.state.put newState
        msgMgr.fifos.state.enq newState

  checkEvalState :: Wire State <- mkWire
  isInCheck :: Wire Bool <- mkWire

  hasMoves :: Reg Bool <- mkReg False

  rules
    "handle_GetState": when GetState <- msgMgr.fifos.command.first ==> do
      eval.state.put state
      msgMgr.fifos.state.enq state
      msgMgr.fifos.command.deq
    "handle_Move": when Move m <- msgMgr.fifos.command.first ==> do
      updateState $ move m state
      msgMgr.fifos.command.deq
    "handle_GetSearchMove": when GetSearchMove <- msgMgr.fifos.command.first ==> do
      searchCore.query.put $ SearchQuery {state=state; depth=searchDepth;}
      msgMgr.fifos.command.deq
    "handle_Reset": when Reset <- msgMgr.fifos.command.first ==> do
      updateState $ initialState
      msgMgr.fifos.command.deq

    -- This is split into seperate rules with wires to avoid excessive compilation times caused by aggressive inlining
    "update_moveState": when True ==>
      checkEvalState :=
        case eval.move.first of
          NextMove m -> move m state
          NoMove -> state
    "update_isInCheck": when True ==>
      isInCheck := inCheck checkEvalState.board state.turn

    "report_NextMove": when NextMove m <- eval.move.first ==> do
      if isInCheck
        then noAction
        else do hasMoves := True
                msgMgr.fifos.moves.enq $ NextMove m
      eval.move.deq
    "report_NoMove": when NoMove <- eval.move.first ==> do
      let outcome :: Outcome =
            case (isInCheck, hasMoves) of
              (False, False) -> Draw
              (False, True) -> NoOutcome
              (True, False) -> CheckMate
              (True, True) -> Check
      msgMgr.fifos.moves.enq NoMove
      msgMgr.fifos.outcome.enq outcome
      hasMoves := False
      eval.move.deq
    "report_search_move": when True ==> do
      result <- searchCore.result.get
      msgMgr.fifos.searchMove.enq result.bestMove

  interface
    txData = enc.byte
    rxData = dec.byte
