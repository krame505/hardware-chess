package Driver where

import Chess
import SearchCore
import GenCMsg
import GenCRepr
import GetPut
import Connectable
import Clocks
import COBS
import CShow

data Command = GetState
             | Move Move
             | GetSearchMove { rid :: RequestId; depth :: Depth; }
             | CancelSearch
             | Reset
  deriving (Bits)

data Outcome = NoOutcome | Check | CheckMate | Draw
  deriving (Bits)

interface ChessMsgs =
  command :: Rx 2 2 Command
  state :: Tx 2 2 State
  outcome :: Tx 2 2 Outcome
  moves :: Tx 64 8 MoveResponse
  searchResult :: Tx 2 2 SearchResult

interface ChessDriver =
  txData :: Get (Bit 8)
  rxData :: Put (Bit 8)

  status :: Bit 8  {-# always_ready, always_enabled #-}

{-# verilog mkChessDriver #-}
mkChessDriver :: Module ChessDriver
mkChessDriver = _mkChessDriver

-- Seperate due to the context
_mkChessDriver :: (GenCMsg ChessMsgs rxBytes txBytes) => Module ChessDriver
_mkChessDriver = module
  writeCMsgDecls "chess" (_ :: ChessMsgs)

  enc :: COBSEncoder txBytes <- mkCOBSEncoder
  dec :: COBSDecoder rxBytes <- mkCOBSDecoder
  msgMgr :: MsgManager ChessMsgs rxBytes txBytes <- mkMsgManager

  dec.msg <-> dropSize msgMgr.rxMsg
  msgMgr.txMsg <-> enc.msg

  state :: Reg State <- mkReg initialState
  eval :: MoveEval <- mkMoveEval

  currentClock <- exposeCurrentClock
  searchCoreReset <- mkReset 1 True currentClock
  searchCore <- changeSpecialWires Nothing (Just searchCoreReset.new_rst) Nothing mkDefaultSearchCore

  let updateState newState = do
        state := newState
        eval.state.put newState
        searchCoreReset.assertReset
        msgMgr.fifos.state.enq newState

  checkEvalState :: Wire State <- mkWire
  isInCheck :: Wire Bool <- mkWire

  hasMoves :: Reg Bool <- mkReg False

  rules
    "handle_GetState": when GetState <- msgMgr.fifos.command.first ==> do
      eval.state.put state
      msgMgr.fifos.state.enq state
      msgMgr.fifos.command.deq
    "handle_Move": when Move m <- msgMgr.fifos.command.first ==> do
      updateState $ move m state
      msgMgr.fifos.command.deq
    "handle_GetSearchMove": when GetSearchMove {rid=rid; depth=depth;} <- msgMgr.fifos.command.first, not searchCoreReset.isAsserted ==> do
      searchCore.query.put $ SearchQuery {rid=rid; state=state; depth=depth;}
      msgMgr.fifos.command.deq
    "handle_CancelSearch": when CancelSearch <- msgMgr.fifos.command.first ==> do
      searchCoreReset.assertReset
      msgMgr.fifos.command.deq
    "handle_Reset": when Reset <- msgMgr.fifos.command.first ==> do
      updateState $ initialState
      msgMgr.fifos.command.deq

    -- This is split into seperate rules with wires to avoid excessive compilation times caused by aggressive inlining
    "update_moveState": when True ==>
      checkEvalState :=
        case eval.move.first of
          NextMove m -> move m state
          NoMove -> state
    "update_isInCheck": when True ==>
      isInCheck := inCheck checkEvalState.board state.turn

    "report_NextMove": when NextMove m <- eval.move.first ==> do
      if isInCheck
        then noAction
        else do hasMoves := True
                msgMgr.fifos.moves.enq $ NextMove m
      eval.move.deq
    "report_NoMove": when NoMove <- eval.move.first ==> do
      let outcome :: Outcome =
            if state.lastProgressMove >= 50 then Draw else
            case (isInCheck, hasMoves) of
              (False, False) -> Draw
              (False, True) -> NoOutcome
              (True, False) -> CheckMate
              (True, True) -> Check
      msgMgr.fifos.moves.enq NoMove
      msgMgr.fifos.outcome.enq outcome
      hasMoves := False
      eval.move.deq
    "report_search_move": when not searchCoreReset.isAsserted ==> do
      result <- searchCore.result.get
      msgMgr.fifos.searchResult.enq result

  interface
    txData = enc.byte
    rxData = dec.byte
    status = searchCore.status
