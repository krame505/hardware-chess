
import "BDPI" function ActionValue#(Int#(32)) rxData();
import "BDPI" function Action txData(Bit#(8) data);
