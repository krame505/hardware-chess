package HwTop where

import Driver
import RS232
import GetPut
import Connectable
import Clocks

interface Top =
  tx :: Bit 1 {-# always_ready, always_enabled #-}
  rx :: Bit 1 -> Action {-# always_ready, always_enabled, prefix="", arg_names = [rx] #-}

clockFreq :: Integer
clockFreq = 100000000

clockDivisor :: Integer
clockDivisor = 2

baud :: Integer
baud = 115200

{-# verilog mkTop #-}
mkTop :: Module Top
mkTop = module
  clockDivider <- mkClockDivider clockDivisor
  reset <- mkReset clockDivisor True clockDivider.slowClock
  driver <- changeSpecialWires (Just clockDivider.slowClock) (Just reset.new_rst) Nothing mkChessDriver
  driverTx <- mkConverter 2 driver.txData
  driverRx <- mkConverter 2 driver.rxData

  uart :: UART 8 <- mkUART 8 NONE STOP_1 (fromInteger $ clockFreq / (baud * 16))
  driverTx <-> uart.rx
  uart.tx <-> driverRx

  interface
    tx = uart.rs232.sout
    rx = uart.rs232.sin
