package SearchCore where

import Chess
import FIFO
import FIFOF
import BRAMFIFO
import GetPut
import Connectable
import Vector
import CShow

type Depth = UInt 8
type Score = Int 8
type MoveCount = UInt 8

moveQueueSize :: Integer
moveQueueSize = 100

pieceValue :: PieceKind -> Score
pieceValue Pawn = 1
pieceValue Knight = 3
pieceValue Bishop = 3
pieceValue Rook = 5
pieceValue Queen = 9
pieceValue King = 0

heuristicScore :: State -> Score
heuristicScore state =
  let squareScore Nothing = 0
      squareScore (Just piece) =
        (if piece.color == state.turn then id else negate) $ pieceValue piece.kind
  in foldr1 (+) $ map squareScore $ concat state.board

struct SearchQuery =
  state :: State
  depth :: Depth
 deriving (Bits)

struct SearchResult =
  bestMove :: Maybe Move
  score :: Score
  depth :: Depth
 deriving (Bits)

interface Frame =
  putState :: State -> Bool -> Action
  putScore :: Score -> ActionValue Bool
  state :: State
  hasMove :: Bool
  score :: Score
  moves :: FIFOF Move

mkFrame :: Module Frame
mkFrame = module
  state <- mkReg _
  inCheck <- mkReg False
  moves <- {- mkSizedBRAMFIFOF -} mkSizedFIFOF moveQueueSize
  hasMove <- mkReg False
  bestScore <- mkReg 0

  interface
    putState s c =
      do state := s
         inCheck := c
         hasMove := False
    putScore s =
      do hasMove := True
         let isBestScore = s > bestScore || not hasMove
         if isBestScore then bestScore := s else noAction
         return isBestScore
    state = state
    hasMove = hasMove
    score =
      if hasMove then bestScore
      else if inCheck then minBound + 1  -- Checkmate
      else 0  -- Draw
    moves = moves

interface (SearchCore :: # -> *) maxDepth =
  query :: Put SearchQuery
  result :: Get SearchResult

  status :: Bit 8 {-# always_ready, always_enabled #-}

mkSearchCore :: (Add 1 n maxDepth) => Module (SearchCore maxDepth)
mkSearchCore = module
  queries :: FIFO SearchQuery <- mkFIFO
  results :: FIFO SearchResult <- mkFIFO

  depth :: Reg Depth <- mkReg 0

  stack :: Vector maxDepth Frame <- replicateM mkFrame
  stackSize :: Reg Depth <- mkReg 0
  let topFrame = select stack (stackSize - 1)
      bottomFrame = stack !! 0

  stateMove :: Wire Move <- mkWire
  state :: Wire State <- mkWire
  stateHeuristicScore :: Wire Score <- mkWire
  currentPlayerInCheck :: Wire Bool <- mkWire
  otherPlayerInCheck :: Wire Bool <- mkWire

  eval :: MoveEval <- mkMoveEval
  movesComplete :: Reg Bool <- mkReg True
  let putState frame = do
        frame.putState state otherPlayerInCheck
        eval.state.put state
        movesComplete := False

  bestMove :: Reg Move <- mkReg _
  currentMove :: Reg Move <- mkReg _

  rules
    "get_query_state": when stackSize == 0 ==> state := queries.first.state
    "get_move_state": when stackSize > 0 ==> state := move stateMove topFrame.state

    "eval_state": when True ==> do
      stateHeuristicScore := heuristicScore state
      currentPlayerInCheck := inCheck state.board topFrame.state.turn
      otherPlayerInCheck := inCheck state.board (otherColor topFrame.state.turn)

  let frameRules frameIndex =
        let nextFrame = if frameIndex < valueOf maxDepth - 1 then stack !! (frameIndex + 1) else _
            currentFrame = stack !! frameIndex
            prevFrame = if frameIndex > 0 then stack !! (frameIndex - 1) else _
        in
          rules
            when stackSize > 0, stackSize - 1 == fromInteger frameIndex
              rules
                ("state_move_" +++ integerToString frameIndex): when True ==> stateMove := currentFrame.moves.first

                ("put_NextMove_" +++ integerToString frameIndex): when not movesComplete, NextMove m <- eval.move.first ==> do
                  -- $display (List.foldr (+++) "" $ List.replicate frameIndex "  ") frameIndex " put_NextMove " (cshow m)
                  currentFrame.moves.enq m
                  eval.move.deq
                ("put_NoMove_" +++ integerToString frameIndex): when not movesComplete, NoMove <- eval.move.first ==> do
                  -- $display (List.foldr (+++) "" $ List.replicate frameIndex "  ") frameIndex " put_NoMove"
                  movesComplete := True
                  eval.move.deq
                ("discard_overflow_state_" +++ integerToString frameIndex): when not movesComplete, not currentPlayerInCheck, fromInteger frameIndex < depth, not currentFrame.moves.notFull ==> do
                  $display (List.foldr (+++) "" $ List.replicate frameIndex "  ") frameIndex " discard_overflow_state " (cshow currentFrame.moves.first)
                  currentFrame.moves.deq

                ("ignore_check_state_" +++ integerToString frameIndex): when currentPlayerInCheck ==> do
                  $display (List.foldr (+++) "" $ List.replicate frameIndex "  ") frameIndex " ignore_check_state " (cshow currentFrame.moves.first)
                  currentFrame.moves.deq

                ("heuristic_state_" +++ integerToString frameIndex): when not currentPlayerInCheck, fromInteger frameIndex >= depth ==> do
                  $display (List.foldr (+++) "" $ List.replicate frameIndex "  ") frameIndex " heuristic_state " (cshow currentFrame.moves.first) " " stateHeuristicScore
                  isBestScore <- currentFrame.putScore $ negate stateHeuristicScore
                  if frameIndex == 0 && isBestScore then bestMove := currentFrame.moves.first else noAction
                  currentFrame.moves.deq

                when movesComplete
                  rules
                    ("push_state_" +++ integerToString frameIndex): when not currentPlayerInCheck, fromInteger frameIndex < depth ==> do
                      $display (List.foldr (+++) "" $ List.replicate frameIndex "  ") frameIndex " push_state " (cshow currentFrame.moves.first) " " stateHeuristicScore
                      putState nextFrame
                      if frameIndex == 0 then currentMove := currentFrame.moves.first else noAction
                      currentFrame.moves.deq
                      stackSize := fromInteger frameIndex + 2

                    ("pop_state_" +++ integerToString frameIndex): when frameIndex > 0, not currentFrame.moves.notEmpty ==> do
                      $display (List.foldr (+++) "" $ List.replicate frameIndex "  ") frameIndex " pop_state " currentFrame.score
                      isBestScore <- prevFrame.putScore $ negate currentFrame.score
                      if frameIndex == 1 && isBestScore then bestMove := currentMove else noAction
                      stackSize := fromInteger frameIndex

  addRules $ foldr1 rJoin ((genWith frameRules) :: Vector maxDepth Rules)

  rules
    when movesComplete
      rules
        "push_query_state": when stackSize == 0 ==> do
          $display stackSize " push_query_state " (cshow queries.first)
          depth := queries.first.depth
          putState bottomFrame
          stackSize := 1
          queries.deq

        "pop_result_state": when stackSize == 1, not bottomFrame.moves.notEmpty ==> do
          let result = SearchResult {
                bestMove = if bottomFrame.hasMove then Just bestMove else Nothing;
                score=bottomFrame.score;
                depth=depth;
               }
          $display "  " stackSize " pop_result_state " (cshow result)
          results.enq result
          stackSize := 0

  interface
    query = toPut queries
    result = toGet results
    status = pack movesComplete ++ pack topFrame.moves.notEmpty ++ pack (depth > 0) ++ pack (impCondOf currentPlayerInCheck) ++ ((truncate $ pack stackSize) :: Bit 4)

{-# verilog mkDefaultSearchCore #-}
mkDefaultSearchCore :: Module (SearchCore 8)
mkDefaultSearchCore = mkSearchCore
