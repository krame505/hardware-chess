package Driver where

import Chess
import SearchCore
import DefaultSearchCores
import GenCMsg
import GenCRepr
import GetPut
import ClientServer
import Connectable
import COBS
import CShow
import FIFO

data Command = GetState
             | Move Move
             | Query { rid :: RequestId; move :: Maybe Move; depth :: Depth; alpha :: Maybe Score; beta :: Maybe Score; getMoves :: Bool }
             | CancelSearch
             | Reset
  deriving (Bits)

struct MoveQuery =
  rid :: RequestId
  depth :: Depth
  alpha :: Maybe Score
  beta :: Maybe Score
  getMoves :: Bool
 deriving (Bits)

interface ChessMsgs =
  command :: Rx 2 2 Command
  state :: Tx 2 2 State
  moves :: Tx 64 8 MoveResponse
  searchResult :: Tx 2 2 SearchResult

interface ChessDriver =
  txData :: Get (Bit 8)
  rxData :: Put (Bit 8)

  status :: Bit 16  {-# always_ready, always_enabled #-}

{-# verilog mkChessDriver #-}
mkChessDriver :: Module ChessDriver
mkChessDriver = _mkChessDriver

-- Seperate due to the context
_mkChessDriver :: (GenCMsg ChessMsgs rxBytes txBytes) => Module ChessDriver
_mkChessDriver = module
  writeCMsgDecls "chess" (_ :: ChessMsgs)

  enc :: COBSEncoder txBytes <- mkCOBSEncoder
  dec :: COBSDecoder rxBytes <- mkCOBSDecoder
  msgMgr :: MsgManager ChessMsgs rxBytes txBytes <- mkMsgManager

  dec.msg <-> dropSize msgMgr.rxMsg
  msgMgr.txMsg <-> enc.msg

  state :: Reg State <- mkReg initialState
  moveUpdate <- mkMoveUpdate
  moveQueries :: FIFO (Maybe MoveQuery) <- mkSizedFIFO 4
  searchCore <- mkParallelSearchCore

  searchCore.moves <-> toPut msgMgr.fifos.moves
  searchCore.server.response <-> toPut msgMgr.fifos.searchResult

  rules
    when not moveUpdate.hasRequest
      rules
        "handle_GetState": when GetState <- msgMgr.fifos.command.first ==> do
          $display "handle_GetState"
          msgMgr.fifos.state.enq state
          msgMgr.fifos.command.deq
        "handle_Move": when Move m <- msgMgr.fifos.command.first ==> do
          $display "handle_Move"
          moveUpdate.enq state m
          moveQueries.enq Nothing
          searchCore.clear
          msgMgr.fifos.command.deq
        "handle_Query": when Query {rid; move; depth; alpha; beta; getMoves;} <- msgMgr.fifos.command.first ==> do
          $display "handle_Query"
          case move of
            Just m -> do
              moveUpdate.enq state m
              moveQueries.enq $ Just $ MoveQuery {rid=rid; depth=depth; alpha=alpha; beta=beta; getMoves=getMoves;}
            Nothing ->
              searchCore.server.request.put $ defaultValue {rid=rid; state=state; depth=depth; alpha=alpha; beta=beta; getMoves=getMoves;}
          msgMgr.fifos.command.deq
        "handle_CancelSearch": when CancelSearch <- msgMgr.fifos.command.first ==> do
          $display "handle_CancelSearch"
          searchCore.clear
          msgMgr.fifos.command.deq
        "handle_Reset": when Reset <- msgMgr.fifos.command.first ==> do
          $display "handle_Reset"
          state := initialState
          searchCore.clear
          msgMgr.fifos.command.deq

    "handle_move_update": when moveUpdate.hasRequest ==> do
      $display "handle_move_update"
      case moveQueries.first of
        Nothing -> state := moveUpdate.nextState
        Just (MoveQuery {rid; depth; alpha; beta; getMoves}) ->
          searchCore.server.request.put $ defaultValue {rid=rid; state=moveUpdate.nextState; depth=depth; alpha=alpha; beta=beta; getMoves=getMoves;}
      moveUpdate.deq
      moveQueries.deq

  interface
    txData = enc.byte
    rxData = dec.byte
    status = searchCore.status
