package SearchCore where

import Chess
import FIFO
import FIFOF
import BRAMFIFO
import GetPut
import Connectable
import Vector
import CShow

type RequestId = UInt 8
type Depth = UInt 8
type Score = Int 8
type MoveCount = UInt 8

minScore :: Score
minScore = minBound + 1  -- We want -minScore = maxScore
maxScore :: Score
maxScore = maxBound

moveQueueSize :: Integer
moveQueueSize = 100

pieceValue :: PieceKind -> Score
pieceValue Pawn = 1
pieceValue Knight = 3
pieceValue Bishop = 3
pieceValue Rook = 5
pieceValue Queen = 9
pieceValue King = 0

heuristicScore :: State -> Score
heuristicScore state =
  let squareScore Nothing = 0
      squareScore (Just piece) =
        (if piece.color == state.turn then id else negate) $ pieceValue piece.kind
  in foldr1 (+) $ map squareScore $ concat state.board

struct SearchQuery =
  rid :: RequestId
  state :: State
  depth :: Depth
 deriving (Bits)

struct SearchResult =
  rid :: RequestId
  bestMove :: Maybe Move
  score :: Score
  depth :: Depth
 deriving (Bits)

interface Frame =
  putState :: State -> Bool -> Score -> Score -> Action
  putScore :: Score -> ActionValue Bool
  state :: State
  hasMove :: Bool
  score :: Score
  alpha :: Score
  beta :: Score
  moves :: FIFOF Move

mkFrame :: Module Frame
mkFrame = module
  state <- mkReg _
  inCheck <- mkReg False
  moves <- {- mkSizedBRAMFIFOF -} mkSizedFIFOF moveQueueSize
  hasMove <- mkReg False
  bestScore <- mkReg 0
  alpha <- mkReg minScore
  beta <- mkReg maxScore

  interface
    putState s c a b =
      do state := s
         inCheck := c
         hasMove := False
         alpha := a
         beta := b
    putScore s =
      do hasMove := True
         let isBestScore = s > bestScore || not hasMove
         if isBestScore then bestScore := s else noAction
         if s > alpha then alpha := s else noAction
         return isBestScore
    state = state
    hasMove = hasMove
    score =
      if hasMove then bestScore
      else if inCheck then minScore  -- Checkmate
      else 0  -- Draw
    alpha = alpha
    beta = beta
    moves = moves

interface (SearchCore :: # -> *) maxDepth =
  query :: Put SearchQuery
  result :: Get SearchResult

  status :: Bit 8 {-# always_ready, always_enabled #-}

mkSearchCore :: (Add 1 n maxDepth) => Module (SearchCore maxDepth)
mkSearchCore = module
  queries :: FIFO SearchQuery <- mkFIFO
  results :: FIFO SearchResult <- mkFIFO

  depth :: Reg Depth <- mkReg 0

  stack :: Vector maxDepth Frame <- replicateM mkFrame
  stackSize :: Reg Depth <- mkReg 0
  let topFrame = select stack (stackSize - 1)
      bottomFrame = stack !! 0

  stateMove :: Wire Move <- mkWire
  state :: Wire State <- mkWire
  stateHeuristicScore :: Wire Score <- mkWire
  currentPlayerInCheck :: Wire Bool <- mkWire
  otherPlayerInCheck :: Wire Bool <- mkWire

  eval :: MoveEval <- mkMoveEval
  movesComplete :: Reg Bool <- mkReg True
  let pushState frame alpha beta = do
        frame.putState state otherPlayerInCheck alpha beta
        eval.state.put state
        movesComplete := False

  bestMove :: Reg Move <- mkReg _
  currentMove :: Reg Move <- mkReg _

  rules
    "get_query_state": when stackSize == 0 ==> state := queries.first.state
    "get_move_state": when stackSize > 0 ==> state := move stateMove topFrame.state

    "eval_state": when True ==> do
      stateHeuristicScore := heuristicScore state
      currentPlayerInCheck := inCheck state.board topFrame.state.turn
      otherPlayerInCheck := inCheck state.board (otherColor topFrame.state.turn)

  let frameRules frameIndex =
        let nextFrame = if frameIndex < valueOf maxDepth - 1 then stack !! (frameIndex + 1) else _
            currentFrame = stack !! frameIndex
            prevFrame = if frameIndex > 0 then stack !! (frameIndex - 1) else _
            isDraw = state.lastProgressMove >= 50
            isTerminal = fromInteger frameIndex >= depth - 1 || isDraw
            depthStr = (List.foldr (+++) "" $ List.replicate (frameIndex + 1) "  ") +++ integerToString (frameIndex + 1)
        in
          rules
            when stackSize > 0, stackSize - 1 == fromInteger frameIndex
              rules
                ("cutoff_" +++ integerToString frameIndex): when frameIndex > 0, currentFrame.alpha >= currentFrame.beta ==> do
                  $display depthStr " cutoff " currentFrame.score
                  prevFrame.putScore $ negate currentFrame.score
                  stackSize := fromInteger frameIndex
                  movesComplete := True
                  currentFrame.moves.clear
                  eval.clear

                when currentFrame.alpha < currentFrame.beta
                  rules
                    ("state_move_" +++ integerToString frameIndex): when True ==> stateMove := currentFrame.moves.first

                    ("put_NextMove_" +++ integerToString frameIndex): when not movesComplete, NextMove m <- eval.move.first ==> do
                      -- $display depthStr " put_NextMove " (cshow m)
                      currentFrame.moves.enq m
                      eval.move.deq
                    ("put_NoMove_" +++ integerToString frameIndex): when not movesComplete, NoMove <- eval.move.first ==> do
                      -- $display depthStr " put_NoMove"
                      movesComplete := True
                      eval.move.deq
                    ("discard_overflow_state_" +++ integerToString frameIndex): when not movesComplete, not currentPlayerInCheck, not isTerminal, not currentFrame.moves.notFull ==> do
                      $display depthStr " discard_overflow_state " (cshow currentFrame.moves.first)
                      currentFrame.moves.deq

                    ("ignore_check_state_" +++ integerToString frameIndex): when currentPlayerInCheck ==> do
                      $display depthStr " ignore_check_state " (cshow currentFrame.moves.first)
                      currentFrame.moves.deq

                    ("heuristic_state_" +++ integerToString frameIndex): when not currentPlayerInCheck, isTerminal ==> do
                      $display depthStr " heuristic_state " (cshow currentFrame.moves.first) " " stateHeuristicScore
                      isBestScore <- currentFrame.putScore $ if isDraw then 0 else negate stateHeuristicScore
                      if frameIndex == 0 && isBestScore then bestMove := currentFrame.moves.first else noAction
                      currentFrame.moves.deq

                    when movesComplete
                      rules
                        ("push_state_" +++ integerToString frameIndex): when not currentPlayerInCheck, not isTerminal ==> do
                          $display depthStr " push_state " (cshow currentFrame.moves.first) " " stateHeuristicScore
                          pushState nextFrame (negate currentFrame.beta) (negate currentFrame.alpha)
                          if frameIndex == 0 then currentMove := currentFrame.moves.first else noAction
                          currentFrame.moves.deq
                          stackSize := fromInteger frameIndex + 2

                        ("pop_state_" +++ integerToString frameIndex): when frameIndex > 0, not currentFrame.moves.notEmpty ==> do
                          $display depthStr " pop_state " currentFrame.score
                          isBestScore <- prevFrame.putScore $ negate currentFrame.score
                          if frameIndex == 1 && isBestScore then bestMove := currentMove else noAction
                          stackSize := fromInteger frameIndex

  addRules $ foldr1 rJoin ((genWith frameRules) :: Vector maxDepth Rules)

  rules
    when movesComplete
      rules
        "invalid_query_depth": when stackSize == 0, queries.first.depth > fromInteger (valueOf maxDepth) ==> do
          $display (0 :: Depth) " invalid_query_depth " (cshow queries.first)
          results.enq $ SearchResult {rid=queries.first.rid; bestMove=Nothing; score=bottomFrame.score; depth=queries.first.depth;}
          queries.deq

        "push_query_state": when stackSize == 0, queries.first.depth <= fromInteger (valueOf maxDepth) ==> do
          $display (0 :: Depth) " push_query_state " (cshow queries.first)
          depth := queries.first.depth
          pushState bottomFrame minScore maxScore
          stackSize := 1

        "pop_result_state": when stackSize == 1, not bottomFrame.moves.notEmpty || bottomFrame.alpha >= bottomFrame.beta ==> do
          let result = SearchResult {
                rid = queries.first.rid;
                bestMove = if bottomFrame.hasMove then Just bestMove else Nothing;
                score = bottomFrame.score;
                depth = depth;
               }
          $display "  " (1 :: Depth) " pop_result_state " (cshow result)
          results.enq result
          queries.deq
          stackSize := 0
          bottomFrame.moves.clear
          eval.clear

  interface
    query = toPut queries
    result = toGet results
    status = ((truncate $ pack depth) :: Bit 4) ++ ((truncate $ pack stackSize) :: Bit 4)

{-# verilog mkDefaultSearchCore #-}
mkDefaultSearchCore :: Module (SearchCore 15)
mkDefaultSearchCore = mkSearchCore
