package VSimTop where

import Chess
import SearchCore
import CShow
import GetPut
import ClientServer

searchDepth :: Depth
searchDepth = 3

{-# verilog sysChessVSim #-}
sysChessVSim :: Module Empty
sysChessVSim = module
  searchCore <- mkParallelSearchCore
  state <- mkReg initialState

  init <- mkReg False
  rules
    "init": when not init ==> do
      $display (cshow state)
      searchCore.server.request.put $ SearchQuery {rid=0; state=state; depth=searchDepth;}
      init := True
    "move": when init ==> do
      result <- searchCore.server.response.get
      $display (cshow result)
      case result.bestMove of
        Just m -> do
          let newState = move m state
          $display newState
          state := newState
          searchCore.server.request.put $ SearchQuery {rid=0; state=newState; depth=searchDepth;}
        Nothing -> $finish
