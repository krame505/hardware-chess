package VSimTop where

import ChessState
import MoveUpdate
import SearchCore
import ShallowSearchCores
import CShow
import GetPut
import ClientServer

searchDepth :: Depth
searchDepth = 3

{-# verilog sysChessVSim #-}
sysChessVSim :: Module Empty
sysChessVSim = module
  searchCore <- mkShallowParallelSearchCore
  moveUpdate <- mkMoveUpdate
  state <- mkReg initialState

  init <- mkReg False
  rules
    "init": when not init ==> do
      $display (cshow state)
      searchCore.server.request.put $ defaultValue {rid=0; state=state; depth=searchDepth;}
      init := True
    "get_result": when init ==> do
      result <- searchCore.server.response.get
      $display (cshow result)
      case result.bestMove of
        Just m -> moveUpdate.enq state m
        Nothing -> $finish
    "put_query": when init ==> do
      $display moveUpdate.nextState
      state := moveUpdate.nextState
      searchCore.server.request.put $ defaultValue {rid=0; state=moveUpdate.nextState; depth=searchDepth;}
      moveUpdate.deq
