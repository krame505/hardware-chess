package DefaultHeuristic where

import Vector
import BuildVector
import Chess
import SearchCore

type ScoreWeight = UInt 4

weightScore :: Score -> ScoreWeight -> Score
weightScore s w = s * zeroExtend (unpack $ pack w)

struct Config =
  materialValue :: ScoreWeight
  centerControlValue :: ScoreWeight
  extendedCenterControlValue :: ScoreWeight
  castleValue :: ScoreWeight
  pawnStructureValue :: ScoreWeight
 deriving (Bits)

instance DefaultValue Config where
  defaultValue =
    interface Config
      materialValue = 5
      centerControlValue = 2
      extendedCenterControlValue = 1
      castleValue = 9
      pawnStructureValue = 1

pieceValue :: PieceKind -> Score
pieceValue Pawn = 1
pieceValue Knight = 3
pieceValue Bishop = 3
pieceValue Rook = 5
pieceValue Queen = 9
pieceValue King = 0

centerPositions :: Vector 4 Position
centerPositions = vec (Position {rank=3; file=3;}) (Position {rank=3; file=4;}) (Position {rank=4; file=3;}) (Position {rank=4; file=4;})

extendedCenterPositions :: Vector 12 Position
extendedCenterPositions = vec
  (Position {rank=2; file=2;}) (Position {rank=2; file=3;}) (Position {rank=2; file=4;}) (Position {rank=2; file=5;})
  (Position {rank=3; file=2;}) (Position {rank=3; file=5;}) (Position {rank=4; file=2;}) (Position {rank=4; file=5;})
  (Position {rank=5; file=2;}) (Position {rank=5; file=3;}) (Position {rank=5; file=4;}) (Position {rank=5; file=5;})

whitePawnPositions :: Vector (TMul 7 8) Position
whitePawnPositions = concat $ genWith (\ rank -> (genWith (\ file -> Position {rank=fromInteger rank; file=fromInteger file;})) :: Vector 8 Position)

blackPawnPositions :: Vector (TMul 7 8) Position
blackPawnPositions = concat $ genWith (\ rank -> (genWith (\ file -> Position {rank=fromInteger rank + 1; file=fromInteger file;})) :: Vector 8 Position)

pawnStructureScore :: Board -> Color -> Position -> Score
pawnStructureScore board turn pos =
  let isTurnPawn p = selectPos board p == Just (Piece {color=turn; kind=Pawn;})
  in
    if isTurnPawn pos
    then
      (if pos.rank > 0 && pos.file > 0 && isTurnPawn (Position {rank=pos.rank - 1; file=pos.file - 1;}) then 1 else 0) +
      (if pos.rank > 0 && pos.file < 7 && isTurnPawn (Position {rank=pos.rank - 1; file=pos.file + 1;}) then 1 else 0) +
      (if pos.file > 0 && isTurnPawn (Position {rank=pos.rank; file=pos.file - 1;}) then negate 1 else 0)
    else 0

defaultHeuristic :: Heuristic Config
defaultHeuristic config state =
  let squareScore :: Maybe Piece -> Score
      squareScore Nothing = 0
      squareScore (Just piece) =
        (if piece.color == state.turn then id else negate) $ pieceValue piece.kind

      controlScore :: ScoreWeight -> Position -> Score
      controlScore score pos =
        let centerThreats = numThreats state.board (otherColor state.turn) pos + (if isOccupied state.board state.turn pos then 1 else 0)
            centerOtherThreats = numThreats state.board state.turn pos + (if isOccupied state.board (otherColor state.turn) pos then 1 else 0)
        in if centerThreats > centerOtherThreats then unpack $ pack $ extend score
           else if centerThreats < centerOtherThreats then negate $ unpack $ pack $ extend score
           else 0

      castleScore = unpack $ pack $ extend config.castleValue
      whitePawnStructureScore = foldr1 (+) $ map (pawnStructureScore state.board White) whitePawnPositions
      blackPawnStructureScore = foldr1 (+) $ map (pawnStructureScore state.board Black) blackPawnPositions

  in (foldr1 (+) $ map squareScore $ concat state.board) `weightScore` config.materialValue +
     (foldr1 (+) $ map (controlScore config.centerControlValue) centerPositions) +
     (foldr1 (+) $ map (controlScore config.extendedCenterControlValue) extendedCenterPositions) +
     (if state.whiteHist.castled then if state.turn == White then castleScore else negate castleScore else 0) +
     (if state.blackHist.castled then if state.turn == Black then castleScore else negate castleScore else 0) +
     (if state.turn == White then id else negate) (whitePawnStructureScore - blackPawnStructureScore) `weightScore` config.pawnStructureValue
