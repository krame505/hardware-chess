package Driver where

import Chess
import GenCMsg
import GenCRepr
import GetPut
import Connectable
import COBS
import CShow

data Command = GetState
             | Reset
  deriving (Bits)

interface ChessMsgs =
  command :: Rx 2 2 Command
  state :: Tx 2 2 State
  moves :: Tx 64 8 MoveResponse

interface ChessDriver =
  txData :: Get (Bit 8)
  rxData :: Put (Bit 8)

mkChessDriver :: (GenCMsg ChessMsgs rxBytes txBytes) => Module ChessDriver
mkChessDriver = module
  writeCMsgDecls "chess" (_ :: ChessMsgs)

  enc :: COBSEncoder txBytes <- mkCOBSEncoder
  dec :: COBSDecoder rxBytes <- mkCOBSDecoder
  msgMgr :: MsgManager ChessMsgs rxBytes txBytes <- mkMsgManager

  dec.msg <-> dropSize msgMgr.rxMsg
  msgMgr.txMsg <-> enc.msg

  state :: Reg State <- mkReg initialState

  eval :: StateEval <- mkStateEval
  eval.moves <-> toPut msgMgr.fifos.moves

  rules
    "handle_command": when True ==> do
      let newState =
            case msgMgr.fifos.command.first of
              GetState -> state
              Reset -> initialState
      state := newState
      eval.state.put newState
      msgMgr.fifos.state.enq newState
      msgMgr.fifos.command.deq

  interface
    txData = enc.byte
    rxData = dec.byte
