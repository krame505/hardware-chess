package HwTop where

import Driver
import RS232
import GetPut
import Connectable

interface Top =
  tx :: Bit 1 {-# always_ready, always_enabled #-}
  rx :: Bit 1 -> Action {-# always_ready, always_enabled, prefix="", arg_names = [rx] #-}

clockFreq :: Integer
clockFreq = 100000000

baud :: Integer
baud = 115200

{-# verilog mkTop #-}
mkTop :: Module Top
mkTop = module
  driver <- mkChessDriver

  uart :: UART 8 <- mkUART 8 NONE STOP_1 (fromInteger $ clockFreq / (baud * 16))
  driver.txData <-> uart.rx
  uart.tx <-> driver.rxData

  interface
    tx = uart.rs232.sout
    rx = uart.rs232.sin
