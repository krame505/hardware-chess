package Driver where

import Chess
import SearchCore
import DefaultSearchCores
import GenCMsg
import GenCRepr
import GetPut
import ClientServer
import Connectable
import COBS
import CShow
import FIFO

data Command = GetState
             | Move Move
             | Query { rid :: RequestId; move :: Maybe Move; depth :: Depth; resetAlpha :: Bool; getMoves :: Bool }
             | CancelSearch
             | Reset
  deriving (Bits)

interface ChessMsgs =
  command :: Rx 2 2 Command
  state :: Tx 2 2 State
  moves :: Tx 64 8 MoveResponse
  searchResult :: Tx 2 2 SearchResult

interface ChessDriver =
  txData :: Get (Bit 8)
  rxData :: Put (Bit 8)

  status :: Bit 16  {-# always_ready, always_enabled #-}

data Task = MoveUpdate
          | MoveQuery { rid :: RequestId; depth :: Depth; resetAlpha :: Bool; getMoves :: Bool }
  deriving (Bits)

{-# verilog mkChessDriver #-}
mkChessDriver :: Module ChessDriver
mkChessDriver = _mkChessDriver

-- Seperate due to the context
_mkChessDriver :: (GenCMsg ChessMsgs rxBytes txBytes) => Module ChessDriver
_mkChessDriver = module
  writeCMsgDecls "chess" (_ :: ChessMsgs)

  enc :: COBSEncoder txBytes <- mkCOBSEncoder
  dec :: COBSDecoder rxBytes <- mkCOBSDecoder
  msgMgr :: MsgManager ChessMsgs rxBytes txBytes <- mkMsgManager

  dec.msg <-> dropSize msgMgr.rxMsg
  msgMgr.txMsg <-> enc.msg

  state :: Reg State <- mkReg initialState
  moveTasks :: FIFO (Move, Task) <- mkSizedFIFO moveQueueSize
  moveUpdate <- mkMoveUpdate
  tasks :: FIFO Task <- mkFIFO
  alpha :: Reg Score <- mkReg minScore
  searchCore <- mkParallelSearchCore

  searchCore.moves <-> toPut msgMgr.fifos.moves

  let clear = do
        moveTasks.clear
        moveUpdate.clear
        tasks.clear
        searchCore.clear

      resultRule =
        rules
          "handle_search_result": when True ==> do
            result <- searchCore.server.response.get
            $display "handle_search_result " (cshow result)
            msgMgr.fifos.searchResult.enq result
            if negate result.score > alpha
              then alpha := negate result.score
              else noAction

      commandRules =
        rules
          "handle_GetState": when GetState <- msgMgr.fifos.command.first ==> do
            $display "handle_GetState"
            msgMgr.fifos.state.enq state
            msgMgr.fifos.command.deq
          "handle_Move": when Move m <- msgMgr.fifos.command.first ==> do
            $display "handle_Move"
            moveTasks.enq (m, MoveUpdate)
            msgMgr.fifos.command.deq
          "handle_direct_Query": when Query {rid; move=Nothing; depth; resetAlpha=_; getMoves;} <- msgMgr.fifos.command.first ==> do
            $display "handle_direct_Query"
            searchCore.server.request.put $ defaultValue {rid=rid; state=state; depth=depth; getMoves=getMoves;}
            msgMgr.fifos.command.deq
          "handle_move_Query": when Query {rid; move=Just m; depth; resetAlpha; getMoves;} <- msgMgr.fifos.command.first ==> do
            $display "handle_Query"
            moveTasks.enq (m, MoveQuery {rid=rid; depth=depth; resetAlpha=resetAlpha; getMoves=getMoves;})
            msgMgr.fifos.command.deq
          "handle_CancelSearch": when CancelSearch <- msgMgr.fifos.command.first ==> do
            $display "handle_CancelSearch"
            clear
            msgMgr.fifos.command.deq
          "handle_Reset": when Reset <- msgMgr.fifos.command.first ==> do
            $display "handle_Reset"
            state := initialState
            clear
            msgMgr.fifos.command.deq

          "put_move_update": when (m, t) <- moveTasks.first ==> do
            $display "put_move_update"
            moveUpdate.enq state m
            tasks.enq t
            moveTasks.deq

      moveUpdateRule =
        rules
          "handle_move_update": when True ==> do
            $display "handle_move_update " (cshow tasks.first)
            case tasks.first of
              MoveUpdate -> do
                state := moveUpdate.nextState
                msgMgr.fifos.state.enq moveUpdate.nextState
              MoveQuery {rid; depth; resetAlpha=False; getMoves} ->
                searchCore.server.request.put $ defaultValue {rid=rid; state=moveUpdate.nextState; depth=depth; beta=Just $ negate alpha; getMoves=getMoves;}
              MoveQuery {rid; depth; resetAlpha=True; getMoves} -> do
                alpha := minScore
                searchCore.server.request.put $ defaultValue {rid=rid; state=moveUpdate.nextState; depth=depth; getMoves=getMoves;}
            moveUpdate.deq
            tasks.deq

  addRules $ resultRule <+ commandRules <+ moveUpdateRule

  interface
    txData = enc.byte
    rxData = dec.byte
    status = searchCore.status
