package SimTop where

import Driver
#ifdef TEST
import TestDriver
#else
import GameDriver
#endif
import GetPut
import PTY

mkDriver :: Module Driver
#ifdef TEST
mkDriver = mkChessTestDriver
#else
mkDriver = mkChessDriver
#endif

{-# verilog sysChessSim #-}
sysChessSim :: Module Empty
sysChessSim = module
  driver <- mkDriver

  -- Wait for first byte to be recieved before sending data
  writeEnable <- mkReg False

  rules
    "tx": when writeEnable ==> do
      c <- driver.txData.get
      txData c

    "rx": when True ==> do
      c <- rxData
      if c /= negate 1
        then do driver.rxData.put $ truncate $ pack c
                writeEnable := True
        else noAction
